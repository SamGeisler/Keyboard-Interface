module ps2_receive()
(
    input clk, reset;
);


endmodule